module  Part1 (A,F);
  output	F;
  input		A;

  not		G1 (F,A);
endmodule