module  Part3 (A,B,F);
  output	F;
  input		A,B;
  
  or		G1 (F,A,B);
endmodule