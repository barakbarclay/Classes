module  Part2 (A,B,F);
  output	F;
  input		A,B;
  
  and		G1 (F,A,B);
endmodule